`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/09/2025 09:38:53 AM
// Design Name: 
// Module Name: exam03_var_module
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module watch(
    input clk, reset_p,
    input [2:0] btn,
    output reg [7:0] sec, min);
    
    reg set_watch; //1이면 set 0이면 watch
    always @(posedge clk, posedge reset_p)begin
        if(reset_p)set_watch = 0;
        else if(btn[0])set_watch = ~set_watch;
    end
    
    integer cnt_sysclk;
    always@(posedge clk, posedge reset_p)begin
        if(reset_p)begin
            cnt_sysclk = 0;
            sec = 0;
            min = 0;
        end
        else begin
            if(set_watch) begin
                if(btn[1])begin
                    if(sec >=59) sec= 0;
                    else sec= sec+1;
                end
                if(btn[2]) begin
                    if(min >=59) min= 0;
                    else min= min+1;
                end
            end
            else begin
                if(cnt_sysclk >= 27'd99_999_999)begin
                    cnt_sysclk = 0;
                    if(sec>=59)begin
                        sec=0;
                        if(min>=59) min= 0;
                        else min=min+1;
                    end
                    else sec = sec+1;
                end
                else cnt_sysclk =cnt_sysclk +1;
            end
        end
    
    end
endmodule

module cook_timer(
    input clk, reset_p,
    input btn_start, inc_sec, inc_min, alarm_off,
    output reg [7:0] sec, min,
    output reg alarm);

    reg dcnt_set;
    reg [7:0] m_sec,m_min;
    always @(posedge clk, posedge reset_p)begin
        if(reset_p)begin
            dcnt_set=0;
            alarm=0;
        end
        else begin
            if(btn_start && !(sec==0 &&min==0))dcnt_set= ~dcnt_set; //
            if(sec ==0 && min ==0 && dcnt_set) begin
                dcnt_set = 0;
                alarm=1;
            end
            if(alarm_off || inc_sec ||inc_min)alarm=0;
            if(alarm_off && !dcnt_set && !(sec==0 &&min==0))begin
                m_min=min;
                m_sec=sec;
            end  
        end
    end
    
    integer cnt_sysclk;
    always @(posedge clk, posedge reset_p)begin
        if(reset_p)begin
            cnt_sysclk= 0;
            sec= 0;
            min= 0;
        end
        else begin
            if(dcnt_set)begin
                if(cnt_sysclk >=99_999_999)begin
                    cnt_sysclk =0;
                    if(sec ==0 && min)begin
                        sec=59;
                        min= min-1;
                    end
                    else sec= sec-1;
                end
                else cnt_sysclk= cnt_sysclk +1;
            end
            else begin
                if(inc_sec)begin
                   if(sec >=59)sec=0;
                   else sec= sec+ 1;
                end
                if(inc_min)begin
                   if(min >=59)min=0;
                   else min= min+ 1;
                end
                if(alarm_off && !dcnt_set && sec ==0 && min ==0 )begin
                    min=m_min;
                    sec=m_sec;
                end
            end
        end
    end
    
endmodule




