`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/17/2025 02:03:06 PM
// Design Name: 
// Module Name: tb_dht11_cntr
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_dht11_cntr();
    
    localparam [7:0] humi_value = 8'd70;
    localparam [7:0] tmpr_value = 8'd25;
    localparam [7:0] check_sum = humi_value + tmpr_value;
    localparam [39:0] data = {humi_value, 8'd0,tmpr_value,8'd0,check_sum};

    reg clk, reset_p;
    tri1 dht11_data;  //pull-up 달린 와이어 임피던스일때 1 시뮬레이션 할때만 사용 
    wire  [7:0] humidity, temperature;
    
    reg dout,wr_e;
    assign dht11_data = wr_e ? dout: 'bz;
    
    dht11_cntr DUT( clk, reset_p, dht11_data,
                       humidity, temperature); 
                       
     initial begin
        clk =0;
        reset_p = 1;
        wr_e = 0;
        dout = 0;
     end
     
     always #5 clk = ~clk;
     
     integer i;
     initial begin
        #10;
        reset_p = 0; #10;
        wait(!dht11_data); // wait 문은 기다린다. 
        wait(dht11_data);  //1이 되기를 기다린다.
        #20_000;
        dout =0; wr_e = 1; #80_000;
        wr_e = 0; #80_000;
        wr_e = 1;
        for (i=0; i<40; i= i+1)begin
            dout= 0; #50_000;
            dout= 1;
            if(data[39-i]) #70_000;
            else #27_000;
        end
        dout= 0; #10;
        wr_e = 0; #1000;
        $stop;
     end
    
    
endmodule
















