`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/09/2025 02:18:49 PM
// Design Name: 
// Module Name: tb_SISO
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
/////////////////////////////////////////////////////////////////////////////////
module tb_SISO();
    
    reg clk, reset_p;
    reg d;
    reg en;
    wire f;
    
    localparam [7:0] data = 8'b1011_1100;  //파라미터는 상수  bc
    
    SISO DUT(.clk(clk), .reset_p(reset_p), .d(d), .en(en), .f(f));

    initial begin
        clk =0;
        reset_p =1;
        en = 0;
    end
    always #5 clk =~clk; 
    
    integer i;
    initial begin
        #10;
        reset_p=0; en=1;
        for(i=0; i<8; i=i+1)begin
            d= data[i];
            #10;
        end
        en=0;
        #50;   //시뮬레이션에서만 쓰는 문법 시스템 명령어  
        en=1; #80
        $stop;
    end
endmodule



module tb_SIPO();
    
    reg clk, reset_p;
    reg d;
    reg rd_en;
    wire [7:0] q;
   
    
    localparam [7:0] data = 8'b1011_1100;  //파라미터는 상수  bc
    
    SIPO DUT(.clk(clk), .reset_p(reset_p), .d(d) ,.rd_en(rd_en), .q(q));

    initial begin
        clk =0;
        reset_p =1;
        d=0;
        rd_en = 0;
    end
    always #5 clk =~clk; 
    
    integer i;
    initial begin
        #10;
        reset_p=0; rd_en=0;
        for(i=0; i<8; i=i+1)begin
            d= data[i];
            #10;
        end
        rd_en=1;
        #5;   //시뮬레이션에서만 쓰는 문법 시스템 명령어  
        rd_en=0; #80
        $stop;
    end
endmodule



module tb_PISO();
    
    reg clk, reset_p;
    reg [7:0] d;
    reg shift_load;
    wire q;
   
    
    localparam [7:0] data = 8'b1011_1100;  //파라미터는 상수  bc
    
    PISO DUT(.clk(clk), .reset_p(reset_p), .d(d) ,.shift_load(shift_load), .q(q));

    initial begin
        clk =0;
        reset_p =1;
        d=0;
        shift_load = 1;
    end
    always #5 clk =~clk; 
    
    integer i;
    initial begin
        #10;
        reset_p=0; shift_load=0;
            d= data;
            #10;
        
        shift_load=1;
        #80;   //시뮬레이션에서만 쓰는 문법 시스템 명령어  
       
        $stop;
    end
endmodule



